ELF          >    P      @       �6          @ 8  @         @       @       @       �      �                                                                                                                                      E      E                                           $      $                   �-      �=      �=      H      P                   �-      �=      �=      �      �                   8      8      8                                   X      X      X      D       D              S�td   8      8      8                             P�td                           4       4              Q�td                                                  R�td   �-      �=      �=      0      0             /lib64/ld-linux-x86-64.so.2              GNU � �                   GNU ��fy����q�����o��         GNU                                 �            �e�m                                                  J                       "                      f                       u                          "                    __libc_start_main __cxa_finalize printf libc.so.6 GLIBC_2.2.5 GLIBC_2.34 _ITM_deregisterTMCloneTable __gmon_start__ _ITM_registerTMCloneTable              )          ui	   3      ���   ?       �=             0      �=             �      @             @      �?                    �?                    �?                    �?                    �?                     @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            H��H��/  H��t��H���         �5�/  �%�/  @ �%�/  h    ������%�/  f�        1�I��^H��H���PTE1�1�H�==  �O/  �f.�     @ H�=�/  H��/  H9�tH�./  H��t	���    ��    H�=a/  H�5Z/  H)�H��H��?H��H�H��tH��.  H��t��fD  ��    ���=/   u+UH�=�.   H��tH�=�.  �)����d�����.  ]� ��    ���w���UH��H�}��VH�E�� < ~FH�E�� <t;H�E�� ����Hc�Hi�]AL�H�� �������)�k�^)ȉЃ�!��H�E��H�E�H�E�� ��u���]�UH��H�� �E�prtr�E�r%u �E�LHb0�E�0fc H�=<0c3_FfH�0CbGbCdbH�E�H�U�f�E�N H�E�H���?���H�E�H���3���H�E�H���'���H�M�H�U�H�E�H��H��  H�Ǹ    ������    ��H��H���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             
Decrypted string: %s%s%s
  ;4       ����    ����   0���P   ����   �����              zR x�      ����"                  zR x�  $      x���     FJw� ?;*3$"       D   p���              \   Q���o    A�Cj     |   �����    A�C�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  0      �             )                            <             �=                           �=                    ���o    �             p             �      
       �                                           �?                                                       @             �       	              ���o           ���o          ���o           ���o           ���o                                                                                                                                   �=                      6              @      GCC: (Debian 14.2.0-8) 14.2.0                               ��                	     |                  ��                     �                    �              3     �              I     @             U     �=              |     0              �     �=              �    ��                    ��                �      !                   ��                �     �=              �                      �     �?              �                                            J     @              (    @              /   <              5                     H    @              U    9      o       c                      r   @                                 �     @              N    P      "       �    @              �    �      �       �   @              �                      �  "                   �                   Scrt1.o __abi_tag crtstuff.c deregister_tm_clones __do_global_dtors_aux completed.0 __do_global_dtors_aux_fini_array_entry frame_dummy __frame_dummy_init_array_entry revme.c __FRAME_END__ _DYNAMIC __GNU_EH_FRAME_HDR _GLOBAL_OFFSET_TABLE_ __libc_start_main@GLIBC_2.34 _ITM_deregisterTMCloneTable _edata _fini printf@GLIBC_2.2.5 __data_start rot47_decrypt __gmon_start__ __dso_handle _IO_stdin_used _end __bss_start main __TMC_END__ _ITM_registerTMCloneTable __cxa_finalize@GLIBC_2.2.5 _init  .symtab .strtab .shstrtab .interp .note.gnu.property .note.gnu.build-id .note.ABI-tag .gnu.hash .dynsym .dynstr .gnu.version .gnu.version_r .rela.dyn .rela.plt .init .plt.got .text .fini .rodata .eh_frame_hdr .eh_frame .init_array .fini_array .dynamic .got.plt .data .bss .comment                                                                                                                           #             8      8                                     6             X      X      $                              I             |      |                                     W   ���o       �      �      $                             a             �      �      �                           i             p      p      �                              q   ���o                                                 ~   ���o                   0                            �             @      @      �                            �      B                                                �                                                         �                                                         �             @      @                                   �             P      P      �                             �             <      <      	                              �                                                           �                             4                              �             X       X       �                              �             �=      �-                                   �             �=      �-                                   �             �=      �-      �                           �             �?      �/      (                             �             �?      �/                                                @      0                                                @      0                                         0               0                                                         80      x                          	                      �3      �                                                   �5                                

GNP�